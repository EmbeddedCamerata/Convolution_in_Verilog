`ifndef __CONFIG_H__
`define __CONFIG_H__

// `define BRAM_MODE

`endif /* __CONFIG_H__ */